module hello_world();

	initial begin
		$display("\n\t Hello World! This is me learning Verilog again from scratch \n");
	end
endmodule
